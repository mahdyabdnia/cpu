module finaltestbench;
clock clk();
testBench tb2();

endmodule
