module AddAlu(inA,inB,out);
input [0:63]inA;
input [0:63]inB;
output [0:63]out;

assign out=inA+inB;

   
endmodule
